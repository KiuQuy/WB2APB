module wb2apb
  ();
endmodule 
